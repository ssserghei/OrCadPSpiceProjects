** Profile: "SCHEMATIC1-ACSweepNoise"  [ D:\YandexDisk\SSS_WorkHome\SSS_OrCad PSpice\004_AcAnalNotchFilt\004_AcAnalNotchFilt-PSpiceFiles\SCHEMATIC1\ACSweepNoise.sim ] 

** Creating circuit file "ACSweepNoise.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100Hz 1Hz 100kHz
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
