** Profile: "SCHEMATIC1-1_Test"  [ D:\GitHub\OrCadPSpiceProjects\014_DenCh7Ex1_StepResolution\014_dench7ex1_stepresolution-pspicefiles\schematic1\1_test.sim ] 

** Creating circuit file "1_Test.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Maxim\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10m 0 {schedule(0,0, 2m,0.05m, 4m,0.01m, 6m,0.005m, 8m,0.001m)} 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
