** Profile: "SCHEMATIC1-AcSweep"  [ d:\github\orcadpspiceprojects\006_ex2notchfilter\006_ex2notchfilter-pspicefiles\schematic1\acsweep.sim ] 

** Creating circuit file "AcSweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Maxim\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 10 10k
.STEP LIN PARAM Rvalue 24k 30k 1k 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
