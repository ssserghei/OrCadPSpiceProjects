** Profile: "SCHEMATIC1-ACSweep"  [ D:\GitHub\OrCadPSpiceProjects\005_ExActiveNotchFilt\005_ExActiveNotchFilt-PSpiceFiles\SCHEMATIC1\ACSweep.sim ] 

** Creating circuit file "ACSweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\Program Files\Cadence\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 10 10k
.STEP LIN PARAM ratio 0.1 0.9 0.1 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
