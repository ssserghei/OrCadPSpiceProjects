** Profile: "SCHEMATIC1-AcSweepNoise"  [ d:\yandexdisk\sss_workhome\sss_orcad pspice\004_acanalnotchfilt\004_acanalnotchfilt-PSpiceFiles\SCHEMATIC1\AcSweepNoise.sim ] 

** Creating circuit file "AcSweepNoise.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\Program Files\Cadence\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 1 0.5kHz
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
