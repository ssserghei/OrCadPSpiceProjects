** Profile: "SCHEMATIC1-AcSweep"  [ D:\YANDEXDISK\SSS_WORKHOME\SSS_ORCAD PSPICE\003_RESISTORNETWORK\005_NOTCHFILTEX2\005_NOTCHFILTEX2-PSpiceFiles\SCHEMATIC1\AcSweep.sim ] 

** Creating circuit file "AcSweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 10 10k
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
